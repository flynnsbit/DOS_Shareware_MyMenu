# Language: Swedish (CP850)

#### This file is part of the FreeDOS HTML Help Viewer
#### and is licensed under its terms.

# Program Usage Screen Strings
1.0:FreeDOS HTML Help Viewer
1.1:Options
1.2:Visa hj�lp om detta
1.3:Visa denna hj�lptext
1.4:Anv�nd monokrom sk�rm
1.5:Anv�nd f�rgschema
1.6:Anv�nder Ascii ist�llet f�r ut�kade teckenkoder
1.7:Ange HELP codepage nnn (annars anv�nds befintlig)
1.8:Avancerat
1.9:Anger s�kv�g f�r hj�lp
1.10:Om ingen fil anges s� anv�nds index.htm 
1.11:L�ser en annan hj�lpfil �n index.htm
1.12:N�r anv�ndaren trycker F1 eller klickar p� "Hj�lp om Hj�lp"
1.13:HELP l�ser denna fil. Default �r help.htm
1.14:Milj�variabler
1.15:Katalog/mapp som inneh�ller hj�lpfilerna
1.16:Ange /M, /A, F1, F2 f�r att g�ra dem till default

#Error Message Strings
2.0:Kunde ej allokera minne
2.1:Ogiltigt argument
2.2:Man kan endast ange ett (1) hj�lptema i taget
2.3:Kan inte anv�nda b�de /f och /m
2.4:Skriv "HELP /?" f�r beskrivning.
2.5:Ingen exakt tr�ff f�r angivet tema
2.6:Hittade ej hj�lp f�r angivet tema
2.7:Internt Fel: storleks�ndring misslyckades
2.8:Kunde ej l�sa komprimerad fil
2.9:Kunde inte �ppna
2.10:Ziparkivet tomt eller felaktigt
2.11:Hittar ej filen. L�ser f�rsta html-fil i ziparkivet
2.12:Kunde ej hitta html-fil i ziparkivet
2.13:Ange en giltig codepage
2.14:Angiven codepage st�ds ej
2.15:Befintliga codepage �r

#Menu Strings
#### HTML Help will truncate strings 3.0 and 3.1
#### if they exceed 14 characters.
3.0:Avsluta
3.1:Help on Help
#### HTML Help will truncate strings 3.2-3.5
#### if they exceed 10 characters.
3.2:Bak�t
3.3:Fram�t
3.4:Inneh�ll
3.5:S�k

#Button Label Strings
#### HTML Help will truncate strings 4.0-4.2
#### if they exceed 8 characters.
4.0:OK
4.1:Avbryt
4.2:Hj�lp

#Status Bar Strings
5.0:Letar hj�lptema...
5.1:Full s�kning sker...
5.2:(tryck ESC f�r att avbryta)...

#Search Box Strings
#### HTML Help will truncate strings:
####    6.0      if it exceeds 35 characters;
####    6.1      if it exceeds 20 characters;
####    6.2-6.5  if they exceed 28 characters;
####    6.6-6.13 if they exceed 35 characters.
6.0:S�k hj�lp
6.1:S�ktext:
6.2:skilj p� gemener/VERSALER
6.3:endast hela ord
6.4:full s�kning
6.5:p� denna sida
#Help on Search:
6.6:Vad S�k g�r
#Lines 6.7-6.9 describe "Search":
6.7:full s�kning:
6.8:S�ker i alla filer
6.9:i inneh�llsf�rteckningen.
#Line 6.10 can be used if you need more room.
6.11:p� denna sida:
6.12:Letar endast i det aktuella
6.13:dokumentet.

#Search Results Strings
7.0:S�kresultat
7.1:S�kte i alla filer
# The following line, 7.2, is used as "Searched [FILENAME]"
7.2:Genoms�kte
# The following line, 7.3, is used as "for: [TEXT]"
7.3:efter
7.4:,Sorry, s�kresultat kan inte genoms�kas.
7.5:ANV�NDAREN AVSLUTADE (med ESC)
7.6:Inga resultat funna
